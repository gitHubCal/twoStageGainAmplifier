** Profile: "SCHEMATIC1-Vout"  [ C:\Users\Calvin\Desktop\Electronics 2\Project 3\project 3-pspicefiles\schematic1\vout.sim ] 

** Creating circuit file "Vout.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../project 3-pspicefiles/project 3.lib" 
* From [PSPICE NETLIST] section of C:\Users\Calvin\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 5m 0 0.01m 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
